`ifndef INC_RNDW_BC_DEC_PKG
`define INC_RNDW_BC_DEC_PKG

package sort_pkg;

parameter M = 6;
parameter N  = 8;
parameter W  = 4;
parameter Q = $clog(W);

endpackage : sort_pkg
`endif

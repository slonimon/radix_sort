`ifndef INC_RNDW_BC_DEC_PKG
`define INC_RNDW_BC_DEC_PKG

package sort_pkg;

parameter M = 64;
parameter N  = 16;
parameter W  = 1;
parameter Q = $clog2(W);

endpackage : sort_pkg
`endif

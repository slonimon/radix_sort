`ifndef INC_RNDW_BC_DEC_PKG
`define INC_RNDW_BC_DEC_PKG

package sort_pkg;

parameter M = 32;
parameter N  = 7;
parameter W  = 32;

endpackage : sort_pkg
`endif
